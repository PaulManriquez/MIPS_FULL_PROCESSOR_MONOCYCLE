module XOR_gate 
(
	output Y, 
	input A, B
);

assign Y = A ^ B;

endmodule
