module AND_gate 
(
	output Y, 
	input A, B
);

assign Y = A & B;

endmodule